`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:32:22 03/28/2017 
// Design Name: 
// Module Name:    IM 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module IM(Pc, InstrOut);

	 input [63:0]Pc;
	 output [31:0] InstrOut;
	
	 reg [7:0] IM [0:255];


	 assign  InstrOut = {IM[0],IM[1],IM[2],IM[3]};


	 initial
	 begin
	 //load1
	 IM[0] = 8'b11111000;//Load1 beginning 
	 IM[1] = 8'b01000010;// register 5 value
	 IM[2] = 8'b00000000;
	 IM[3] = 8'b00000101;//load1 ending 
	 
	 //load2
	 IM[4] = 8'b11111000;//load2 beginning
	 IM[5] = 8'b01000101;//register 6 value
	 IM[6] = 8'b00000000;
	 IM[7] = 8'b00001010;//load1 ending 
	 
	 //AluOp1
	 
	 //add
	 IM[8] = 8'b10001011;	
	 IM[9] = 8'b00001010;	//add reg5 with reg6 to reg 1
	 IM[10] = 8'b00000000;
	 IM[11] = 8'b10100001;	
	 
	 //subtract
	 IM[12] = 8'b11001011;	
	 IM[13] = 8'b00001010;	//subtract reg5 with reg6 to reg 2
	 IM[14] = 8'b00000000;
	 IM[15] = 8'b10100010;	
	 
	 //and
	 
	 IM[16] = 8'b10001010;	
	 IM[17] = 8'b00001010;	//and reg5 with reg6 to reg 3
	 IM[18] = 8'b00000000;
	 IM[19] = 8'b10100011;
	 
	 //or
	 IM[20] = 8'b10101010;	
	 IM[21] = 8'b00001010;	//or reg5 with reg6 to reg 3
	 IM[22] = 8'b00000000;
	 IM[23] = 8'b10100100;
	 
	 //store
	 
	  //Store 1
	 IM[20] = 8'b11111000;	
	 IM[21] = 8'b00000000;	//Store x1 to 0
	 IM[22] = 8'b10000000;
	 IM[23] = 8'b00000001;
	 
	   //Store 2
	 IM[20] = 8'b11111000;	
	 IM[21] = 8'b00000001;	//Store x2 to 8
	 IM[22] = 8'b00000000;
	 IM[23] = 8'b00000010;
	 
	   //Store 3
	 IM[20] = 8'b11111000;	
	 IM[21] = 8'b00000010;	//Store x3 to 16 
	 IM[22] = 8'b00000000;
	 IM[23] = 8'b00000011;
	 
	   //Store 4
	 IM[20] = 8'b11111000;	
	 IM[21] = 8'b00000100;	//Store x4 to 24
	 IM[22] = 8'b00000000;
	 IM[23] = 8'b00000100;
	 
	
	 end
endmodule
