`timescale 1ns / 1ps


module Adder_Branch(A, B, out);//is to get the sum of PC and Offset
	
	input [63:0]  A;
	input [44:0] B;
	output reg out;
	

endmodule
